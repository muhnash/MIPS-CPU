module Test();
	wire clock;
	wire w1 , w2 ,w3;
	wire out , ZERO;
	reg in1[31:0] , in2[31:0] , alu_control[3:0];
	reg x;
	
	//in1=32'b0000_0000_0000_0000_0000_0000_0000_0000;
	always@(clock) begin 
	x=0;
	in1=32'b00000000000000000000000000000000;
		
		//ALU(in1,in2,alu_control,out,ZERO);
		
		
		
		
		
	end
	
	
	
endmodule
