module MIPS();
/*
[CSE311 Final Project]
[Main Module]
	
#1 ) Single cycle Implementation: (Lecture 1 > slide #20)
=========================================================
	Instruction Set Supported:
	==========================
		� Arithmetic: add, addi	  
		� Load/Store: lw, sw
		� Logic: sll, and, andi, nor
		� Control flow: beq, jal, jr
		� Comparison: slt

*/

endmodule