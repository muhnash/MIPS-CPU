module ShiftLeft_2(out, in);
input in;
output out;

assign out=in<<2;

endmodule