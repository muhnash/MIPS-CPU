module ALUcontrol(out , func , ALUop);
	input func[5:0], ALUop[2:0]; 
	output out; 
	
endmodule 